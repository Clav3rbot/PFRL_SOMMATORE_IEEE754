
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

entity IEEE754_ADDER is
end IEEE754_ADDER;

architecture Behavioral of IEEE754_ADDER is

begin


end Behavioral;

