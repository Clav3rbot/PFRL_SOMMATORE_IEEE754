
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

entity COMPLEMENT2 is
end COMPLEMENT2;

architecture STRUCT of COMPLEMENT2 is

begin


end STRUCT;

