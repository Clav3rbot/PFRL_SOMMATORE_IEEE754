
LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;

ENTITY CONDITIONAL_C2 IS
	GENERIC (M : NATURAL := 8);
	PORT (
		X : IN STD_LOGIC_VECTOR(M - 1 DOWNTO 0);
		S : IN STD_LOGIC;
		Z : OUT STD_LOGIC_VECTOR(M - 1 DOWNTO 0);
		COUT : OUT STD_LOGIC
	);
END CONDITIONAL_C2;

ARCHITECTURE STRUCT OF CONDITIONAL_C2 IS

	COMPONENT CARRY_ADDER IS
		GENERIC (N : NATURAL := M);
		PORT (
			X : IN STD_LOGIC_VECTOR(M - 1 DOWNTO 0);
			CIN : IN STD_LOGIC;
			S : OUT STD_LOGIC_VECTOR(M - 1 DOWNTO 0);
			COUT : OUT STD_LOGIC
		);
	END COMPONENT;

	SIGNAL XXorS : STD_LOGIC_VECTOR(M - 1 DOWNTO 0);
	SIGNAL SExpander : STD_LOGIC_VECTOR(M - 1 DOWNTO 0);
BEGIN
	SExpander <= (OTHERS => S);
	XXorS <= X XOR SExpander;

	U1 : CARRY_ADDER PORT MAP(
		X => XXorS,
		CIN => S,
		S => Z,
		COUT => COUT
	);
END STRUCT;