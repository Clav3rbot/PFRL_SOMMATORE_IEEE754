
LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;

ENTITY SUM IS
	PORT (
		XSIGN : IN STD_LOGIC;
		YSIGN : IN STD_LOGIC;
		XMAN : IN STD_LOGIC_VECTOR (23 DOWNTO 0);
		YMAN : IN STD_LOGIC_VECTOR (23 DOWNTO 0);
		ZMANT : OUT STD_LOGIC_VECTOR(23 DOWNTO 0);
		EXPINCR : OUT STD_LOGIC
	);
END SUM;

ARCHITECTURE RTL OF SUM IS

	COMPONENT CONDITIONAL_C2 IS
		GENERIC (N : NATURAL);
		PORT (
			X : IN STD_LOGIC_VECTOR(N - 1 DOWNTO 0);
			S : IN STD_LOGIC;
			Z : OUT STD_LOGIC_VECTOR(N - 1 DOWNTO 0);
			COUT : OUT STD_LOGIC
		);
	END COMPONENT;

	COMPONENT RIPPLE_CARRY_ADDER IS
		GENERIC (N : NATURAL);
		PORT (
			X : IN STD_LOGIC_VECTOR (N - 1 DOWNTO 0);
			Y : IN STD_LOGIC_VECTOR (N - 1 DOWNTO 0);
			CIN : IN STD_LOGIC;
			S : OUT STD_LOGIC_VECTOR (N - 1 DOWNTO 0);
			COUT : OUT STD_LOGIC
		);
	END COMPONENT;

	SIGNAL OperationLogic : STD_LOGIC;
	SIGNAL C2Mant : STD_LOGIC_VECTOR(23 DOWNTO 0);

BEGIN

	OperationLogic <= XSIGN xor YSIGN;
	
	U1: CONDITIONAL_C2
		generic map(N => 24)
		port map(
			X => YMAN,
			S => OperationLogic,
			Z => C2Mant
		);
		
	U2: RIPPLE_CARRY_ADDER
		generic map(N => 24)
		port map(
			X => XMAN,
			Y => C2Mant,
			CIN => '0',
			S => ZMant,
			COUT => ExpIncr -- importante ! se = 1 => bisogna incrementare l'esponente
		);

END RTL;