LIBRARY ieee;
USE ieee.std_logic_1164.ALL;
ENTITY TB_ADDER_PIPELINE IS
END TB_ADDER_PIPELINE;

ARCHITECTURE behavior OF TB_ADDER_PIPELINE IS
	-- Component Declaration for the Unit Under Test (UUT)

	COMPONENT IEEE754_ADDER
		PORT (
			X : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
			Y : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
			OP : IN STD_LOGIC;
			Z : OUT STD_LOGIC_VECTOR(31 DOWNTO 0);

			CLK : IN STD_LOGIC;
			RST : IN STD_LOGIC
		);
	END COMPONENT;
	--Inputs
	SIGNAL X : STD_LOGIC_VECTOR(31 DOWNTO 0);
	SIGNAL Y : STD_LOGIC_VECTOR(31 DOWNTO 0);
	SIGNAL OP : STD_LOGIC;

	--Service
	SIGNAL RST : STD_LOGIC;
	SIGNAL CLK : STD_LOGIC;

	--Outputs
	SIGNAL Z : STD_LOGIC_VECTOR(31 DOWNTO 0);

	CONSTANT Clk_Period : TIME := 40 ns;
BEGIN

	-- Instantiate the Unit Under Test (UUT)
	uut : IEEE754_ADDER PORT MAP(
		X => X,
		Y => Y,
		OP => OP,
		Z => Z,

		RST => RST,
		CLK => CLK
	);

	CLK_process : PROCESS
	
	BEGIN
		CLK <= '0';
		WAIT FOR Clk_Period/2;
		CLK <= '1';
		WAIT FOR Clk_Period/2;
	END PROCESS;
	
	-- Stimulus process
	PROCESS
	BEGIN
		
		RST <= '1';
		
		WAIT FOR Clk_Period;
		
		RST <= '0';

      -- ordinary numbers
		X <= "01000100101111100011011110101110"; -- 1521.739990234375
		Y <= "01000100101001101010010011001101"; -- 1333.1500244140625
		OP <= '0';

		-- expected output: 01000101001100100110111000111110 - 2854.89013671875 <
		WAIT FOR Clk_Period;
		X <= "00010000100000000000000000000001"; -- 5.048 10E-29
		Y <= "00010000100000000000000000000000"; -- 5.048 10E-29
		OP <= '0';

		-- expected output: 00010001000000000000000000000000 - 1.009742E-28 <
		WAIT FOR Clk_Period;
		X <= "11000001000000010011101101100100"; -- -8.077   
		Y <= "11000001011001100101101000011101"; -- -14.397
		OP <= '1';

		-- expected output: 01000000110010100011110101110010 - 6.3200006 <
		WAIT FOR Clk_Period;
		X <= "01000100101001101010010011001101"; -- 1333.1500244140625
		Y <= "01000100101111100011011110101110"; -- 1521.739990234375  
		OP <= '0';

		-- expected output: 01000101001100100110111000111110 - 2854.8901 <
		WAIT FOR Clk_Period;
		X <= "00010010100000000000000000000001"; -- 8.077E-28  
		Y <= "00010000100000000000000000000000"; -- 5.048E-29
		OP <= '1';

		-- expected output: 00010010011100000000000000000010 - 7.5730657E-28 <

		WAIT FOR Clk_Period;
		X <= "11000001011001100101101000011101"; -- -14.397  
		Y <= "11000001000000010011101101100100"; -- -8.077
		OP <= '0';

		-- expected output: 11000001101100111100101011000000 - -22.473999 <
		WAIT FOR Clk_Period;

		X <= "00010000100000000000000000000001"; -- 5.0487104E-29
		Y <= "00000000100000000000000000000001"; -- 1.1754945E-38
		OP <= '0';
		-- expected output: 00010000100000000000000000000001 - 5.0487104E-29 <

		-- inf
		WAIT FOR Clk_Period;
		X <= "00000000101101100000001010000001"; -- 1.6714959E-38
		Y <= "00000000101101100000001010000000"; -- 1.6714957E-38
		OP <= '1';
		-- expected output: 00000000000000000000000000000001 - 1E-45 < (rounded to zero?)

		WAIT FOR Clk_Period;
		X <= "01000100101111100011011110101110"; -- 1521.739990234375
		Y <= "01000100101111100011011110101110"; -- 1521.739990234375
		OP <= '1';
		-- expected output: 00000000000000000000000000000000 - 0 <

		WAIT FOR Clk_Period;

		X <= "00000011000000000000000001110000"; -- 3.76163214517E-37
		Y <= "00000011000000000000000011110000"; -- 3.76168954235E-37
		OP <= '1';
		-- expected output: 10000000000000000001000000000000 - -5.74E-42 <

		WAIT FOR Clk_Period;

		X <= "10000000011111111111111111111100"; -- -1.1754938E-38
		Y <= "00000000010000000000011000001101"; --  5.879642E-39
		OP <= '0';
		-- expected output : 10000000001111111111100111101111 - -5.875296E-39 <
		
		-- sup
		WAIT FOR Clk_Period;

		X <= "10000000000000000000000000000011"; -- -4E-45
		Y <= "11111111011111111111111111111111"; -- almost infinity
		OP <= '0';
		-- expected output: 11111111011111111111111111111111 - -3.4028235E38 <
		
		WAIT FOR Clk_Period;
		
		X <= "01111111011111111111111111111100"; -- Big numb
		Y <= "01111111000000000000011000001101"; -- Big numb
		OP <= '0';
		-- expected output: 01111111100000000000000000000000 - +inf ?
		-- non va questo ora
		-- non si vede proprio
		
		-- special cases
		WAIT FOR Clk_Period;

		X <= "01111111100000000000000000000000"; -- +inf
		Y <= "01111111100000000000000000000000"; -- +inf
		OP <= '1';
		-- expected output: 01111111111111111111111111111111 - NAN <

		WAIT FOR Clk_Period;

		X <= "11111111100000000000000000000000"; -- -inf
		Y <= "01111111100000000000000000000000"; -- +inf
		OP <= '0';
		-- expected output: 01111111111111111111111111111111 - NAN <

		WAIT FOR Clk_Period;

		X <= "11111111100000000000000000000000"; -- -inf
		Y <= "11111111100000000000000000000000"; -- -inf
		OP <= '0';
		-- expected output: 11111111100000000000000000000000 - -inf <

		WAIT FOR Clk_Period;

		X <= "11111111100000000000000000000000"; -- -inf
		Y <= "11001001100101101011010000111000"; -- -1234567
		OP <= '0';
		-- expected output: 11111111100000000000000000000000 - -inf <

		WAIT FOR Clk_Period; -- +inf - num

		X <= "01111111100000000000000000000000"; -- +inf
		Y <= "11001001100101101011010000111000"; -- -1234567
		OP <= '0';
		-- expected output: 01111111100000000000000000000000 - +inf <

		WAIT FOR Clk_Period; -- inf + 0

		X <= "01111111100000000000000000000000"; -- +inf
		Y <= "00000000000000000000000000000000"; -- 0
		OP <= '0';
		-- expected output: 01111111100000000000000000000000 - +inf <

		WAIT FOR Clk_Period;

		X <= "11111111100000000000000110000000"; -- NAN
		Y <= "11001001100101101011010000111000"; -- -1234567
		OP <= '1';
		-- expected output: 01111111111111111111111111111111 - NAN <

		WAIT FOR Clk_Period;
		
		X <= "01111111100101101011010000111000"; -- NaN
		Y <= "00000000000000000000000000000000"; -- 0
		OP <= '0';
		-- expected output: 01111111111111111111111111111111 - NAN <

		WAIT FOR Clk_Period;

		X <= "01111111100101101011000111101000"; -- NaN
		Y <= "01111111100000000000000000000000"; -- inf
		OP <= '0';
		-- expected output: 01111111111111111111111111111111 - NAN <
		
		WAIT;
	END PROCESS;

END;