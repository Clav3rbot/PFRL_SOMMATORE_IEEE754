
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

entity POST_SUM is
port (
		XCASE : in STD_LOGIC_VECTOR(2 downto 0);
		YCASE : in STD_LOGIC_VECTOR(2 downto 0);
		Z : out STD_LOGIC_VECTOR(31 downto 0)
	);
end POST_SUM;

architecture RTL of POST_SUM is
begin


end RTL;

