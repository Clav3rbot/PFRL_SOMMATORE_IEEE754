LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;

ENTITY NORMALIZER IS
	PORT (
		EXP : IN STD_LOGIC_VECTOR(7 DOWNTO 0);
		MAN : IN STD_LOGIC_VECTOR(26 DOWNTO 0);
		NEXP : OUT STD_LOGIC_VECTOR(7 DOWNTO 0);
		NMAN : OUT STD_LOGIC_VECTOR(25 DOWNTO 0)
	);
END NORMALIZER;

ARCHITECTURE RTL OF NORMALIZER IS

	-- Ci dice la posizione dell'1 più significativo
	COMPONENT PRIORITY_ENCODER
		PORT (
			X : IN STD_LOGIC_VECTOR(26 DOWNTO 0);
			SHIFT : OUT STD_LOGIC_VECTOR(7 DOWNTO 0)
		);
	END COMPONENT;
	
	-- Shifter a sinistra di tante posizioni quanto l'output del modulo PRIORITY_ENCODER
	COMPONENT LEFT_SHIFTER
		PORT (
			X : IN STD_LOGIC_VECTOR(26 DOWNTO 0);
			S : IN STD_LOGIC_VECTOR(7 DOWNTO 0);
			Y : OUT STD_LOGIC_VECTOR(25 DOWNTO 0)
		);
	END COMPONENT;

	-- Decrementare l'esponente
	COMPONENT RIPPLE_CARRY_ADDER

		GENERIC (N : NATURAL);

		PORT (
			X : IN STD_LOGIC_VECTOR (N - 1 DOWNTO 0);
			Y : IN STD_LOGIC_VECTOR (N - 1 DOWNTO 0);
			CIN : IN STD_LOGIC;
			S : OUT STD_LOGIC_VECTOR (N - 1 DOWNTO 0);
			COUT : OUT STD_LOGIC

		);
	END COMPONENT;
	
	COMPONENT MULTIPLEXER_N IS
		GENERIC(N : NATURAL);
		PORT (
        X : IN STD_LOGIC_VECTOR(N - 1 DOWNTO 0);
        Y : IN STD_LOGIC_VECTOR(N - 1 DOWNTO 0);
        S : IN STD_LOGIC;
        Z : OUT STD_LOGIC_VECTOR(N - 1 DOWNTO 0)
    );
	END COMPONENT;	

	SIGNAL ShiftPos : STD_LOGIC_VECTOR(7 DOWNTO 0);
	SIGNAL ManShift : STD_LOGIC_VECTOR(25 DOWNTO 0);
	SIGNAL ExpShift : STD_LOGIC_VECTOR(7 DOWNTO 0);
	SIGNAL NotShiftPos : STD_LOGIC_VECTOR(7 DOWNTO 0);
	SIGNAL AllZero : STD_LOGIC;

BEGIN
	U1 : PRIORITY_ENCODER
	PORT MAP(
		X => MAN,
		SHIFT => ShiftPos
	);

	U2 : LEFT_SHIFTER
	PORT MAP(
		X => MAN,
		S => ShiftPos,
		Y => ManShift
	);
	
	NotShiftPos <= not ShiftPos;
	
	U3 : RIPPLE_CARRY_ADDER
	GENERIC MAP(
		N => 9
	)
	PORT MAP(
		X => '0' & EXP,
		Y => '1' & NotShiftPos,
		CIN => '1',
		S(7 downto 0) => ExpShift,
		S(8) => AllZero
	);
	
	U4: MULTIPLEXER_N
	GENERIC MAP(N => 8)
	PORT MAP(
		X => ExpShift,
		Y => (others => '0'),
		S => AllZero,
		Z => NEXP
	);
	
	U5: MULTIPLEXER_N
	GENERIC MAP(N => 26)
	PORT MAP(
		X => ManShift,
		Y => (others => '0'),
		S => AllZero,
		Z => NMAN
	);

END RTL;
