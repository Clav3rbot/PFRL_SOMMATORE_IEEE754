
LIBRARY ieee;
USE ieee.std_logic_1164.ALL;
USE ieee.numeric_std.ALL;

ENTITY TB_PRE_SUM IS
END TB_PRE_SUM;

ARCHITECTURE behavior OF TB_PRE_SUM IS

	-- Component Declaration
	COMPONENT PRE_SUM
		PORT (
			X : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
			Y : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
			OP : IN STD_LOGIC;
			XSIGN : OUT STD_LOGIC;
			YSIGN : OUT STD_LOGIC;
			XEXP : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
			XMAN : OUT STD_LOGIC_VECTOR (26 DOWNTO 0);
			YMAN : OUT STD_LOGIC_VECTOR (26 DOWNTO 0);
			SPECIAL : OUT STD_LOGIC;
			SPECIAL_RESULT : OUT STD_LOGIC_VECTOR(31 DOWNTO 0)
		);
	END COMPONENT;

	--Inputs
	SIGNAL X : STD_LOGIC_VECTOR(31 DOWNTO 0);
	SIGNAL Y : STD_LOGIC_VECTOR(31 DOWNTO 0);
	SIGNAL op : STD_LOGIC;

	--Outputs
	SIGNAL XSIGN : STD_LOGIC;
	SIGNAL YSIGN : STD_LOGIC;
	SIGNAL XEXP : STD_LOGIC_VECTOR(7 DOWNTO 0);
	SIGNAL XMAN : STD_LOGIC_VECTOR(26 DOWNTO 0);
	SIGNAL YMAN : STD_LOGIC_VECTOR(26 DOWNTO 0);
	SIGNAL SPECIAL : STD_LOGIC;
	SIGNAL SPECIAL_RESULT : STD_LOGIC_VECTOR(31 DOWNTO 0);

BEGIN

	-- Component Instantiation
	uut : PRE_SUM PORT MAP(
		X => X,
		Y => Y,
		OP => OP,
		XSIGN => XSIGN,
		YSIGN => YSIGN,
		XEXP => XEXP,
		XMAN => XMAN,
		YMAN => YMAN,
		SPECIAL => SPECIAL,
		SPECIAL_RESULT => SPECIAL_RESULT
	);

	-- Stimulus process
	stim_proc : PROCESS
	BEGIN
	
		X <= "00000000000000000000000000000000";
		Y <= "00000000000000000000000000000000";
		op <= '0';
		
		WAIT FOR 100 ns;
		
		X <= "10000000000000000000000000000011"; 
		Y <= "11111111011111111111111111111111"; -- almost infinity
		op <= '0';
		
		WAIT FOR 40 ns;
		
		X <= "01000100101111100011011110101110"; -- 1521.739990234375
		Y <= "01000100101111100011011110101110"; -- 1521.739990234375
		op <= '1';
		WAIT FOR 40 ns;
		
		X <= "01000001111010001100110011000000";
		Y <= "01000001111010001100110011000001";
		op <= '0';
		WAIT FOR 40 ns;
		
		X <= "01000001111010001100110011000000";
		Y <= "11000001111010001100110011000000";
		op <= '0';
		WAIT FOR 40 ns;
		
		X <= "01000001111010001100110011000000";
		Y <= "11000001111010001100110011000000";
		op <= '1';
		WAIT FOR 40 ns;
		
		X <= "01000001111010001100110011000000";
		Y <= "11111111111010001100110011000000";
		op <= '1';
		WAIT FOR 40 ns;
		
		X <= "01000001111010001100110011000000";
		Y <= "11111111111010001100110011000000";
		op <= '1';
		WAIT FOR 40 ns;
		
		X <= "00010000100000000000000000000001";
		Y <= "00000000000000000000000000000010";
		op <= '0';
		WAIT FOR 40 ns;
		
		X <= "01111111011111111111111111111111";
		Y <= "00000000000000000000000000000011";
		op <= '0';
		WAIT FOR 40 ns;
		
		X <= "00000000100000000000000000011111";
		Y <= "00000000100000000000000000010001";
		op <= '1';
		WAIT FOR 40 ns;
		
		X <= "00000000011111111111111111111111";
		Y <= "00000000011111111111111111111111";
		op <= '0';
		WAIT FOR 40 ns;
		
		X <= "00010010100000000000000000000001";
		Y <= "00010000100000000000000000000000";
		op <= '1';
		WAIT FOR 40 ns;
		
		X <= "00000011000000000000000001110000";
		Y <= "00000011000000000000000011111000";
		op <= '1';
		WAIT FOR 40 ns;
		
		X <= "01111111100000000000000000000000";
		Y <= "01111111100000000000000000000000";
		op <= '1';
		WAIT FOR 40 ns;
		
		X <= "00000000011111111111111111111111";
		Y <= "00000000011111111111111111111111";
		op <= '0';
		WAIT FOR 40 ns;
		
		X <= "00000000011111111111111111111111";
		Y <= "10000000011111111111111111111111";
		op <= '1';
		WAIT FOR 40 ns;
		
		X <= "10000000000000000000000000000011";
		Y <= "11111111011111111111111111111111";
		op <= '0';
		WAIT FOR 40 ns;
		
		X <= "01111111011111111111111111111111";
		Y <= "01111110000000000000000000000011";
		op <= '0';
		WAIT FOR 40 ns;
		
		X <= "01000100101111100011011110101110";
		Y <= "01000100101001101010010011001101";
		op <= '0';

		WAIT;
	END PROCESS;

END;